* /home/santhosh.ldc20/eSim-Workspace/test_adcBridge/test_adcBridge.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 11:48:45 AM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Vin Net-_U2-Pad2_ adc_bridge_1		
v1  Vin GND pulse		
U1  Vin plot_v1		
U3  Vout plot_v1		
U4  Net-_U2-Pad2_ Vout dac_bridge_1		

.end
