module santhosh_inv(y,a);
	output y;
	input a;
	
	assign y=~a;
	
endmodule
