module santh_inverter(y,a);
	output y;
	input a;
	
	assign y=~a;
	
endmodule
