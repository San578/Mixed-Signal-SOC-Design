* /home/santhosh.ldc20/eSim-Workspace/DFF/DFF.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 09:41:15 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v2  En GND pulse		
v1  in GND pulse		
v3  Net-_SC1-Pad3_ GND DC		
U2  out plot_v1		
U1  in plot_v1		
scmode1  SKY130mode		
SC1  Int_Out Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC2  Int_Out Net-_SC1-Pad2_ Net-_SC2-Pad3_ GND sky130_fd_pr__nfet_01v8		
SC3  Net-_SC2-Pad3_ En GND GND sky130_fd_pr__nfet_01v8		
U4  En plot_v1		
U6  Net-_U3-Pad2_ Net-_SC1-Pad2_ dac_bridge_1		
U5  in Net-_U3-Pad1_ adc_bridge_1		
U12  Int_Out plot_v1		
SC4  Int_Out GND sky130_fd_pr__cap_mim_m3_1		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ santh_inverter		
U8  Int_Out Net-_U7-Pad1_ adc_bridge_1		
U7  Net-_U7-Pad1_ Net-_U7-Pad2_ santh_transmission		
U9  Net-_U7-Pad2_ out dac_bridge_1		

.end
