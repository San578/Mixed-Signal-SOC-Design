module santh_transmission(y,a);
	output y;
	input a;
	
	assign y=a;
	
endmodule
